LAB-3-EXAMPLE-1.cir
R1	1	3	5
R2	2	3	5
R3	2	0	10
R4	4	3	20
R5	3	5	10
V1 1	0	DC	0V
I1	0	4	DC 0A
G1	0	3	2	0	2
IL	0	5	DC	1A
.DC	V1	0	0	1
.PRINT	DC	V(5,0)
.END
