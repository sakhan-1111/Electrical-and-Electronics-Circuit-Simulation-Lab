HOMEWORK_PROBLEM_1.CIR
Is	3	0	DC 0.136092A
R4	1	0	300
R5	2	0	250
R3	1	2	100
R1	3	1	150
R2	3	2	50
.DC	Is	0.136092	0.136092	1
.PRINT	DC	V(1,2)	I(R3)
.END
