LAB-3-EXERCISE-2-NETLIST-3.CIR
R1	1	2	1
R2	2	3	4
R3	3	0	5
R4	3	7	5
R5	6	0	4.8
V1	4	7	DC	0V
Vs	4	2	DC	100V
E1	4	5	2	3	3
F1	1	0	V1	4
RL	5	6	{R}
.PARAM R=10
.DC	PARAM	R	1	20	1
.PROBE
.END

