LAB_2_EXERCISE_3.CIR
R1	1	5	10
R2	1	3	10
R3	1	2	5
R4	2	4	5
R5	2	6	10
V1	5	0	DC 100V
V2	6	0	DC 0V
G1	3	0	1	2	10
H1	4	0	V2	10
.DC	V1	100	100	1
.PRINT DC	V(1) V(2) V(1,2)	I(R5)
.END
