EXANPLE-2-NETLIST.CIR
R1	0 1  1k 
I1	0 1 DC 10mA
C1	0 1  10uF IC=5
.TRAN	20us	150ms	0ms	10us UIC
.PROBE
.END
