test 1.cir
I1         0 1 DC 10A  
R1         1 3  2  
R4         0 3  6  
R2         1 2  3
V1		2	5  DC	0V
F1    3	2	V1	4
R3         0 5  4  
.dc I1	10	10	1
.PRINT DC V(1)V(2)V(3)
.END
