Lab-5-Exercise-1-Netlist.cir
V1	1	0	DC	0	AC	0	SIN	0	100V	60Hz	0	0	0
C1	3	0	10uF
R1	1	2	31.25
R2	1	3	30
L1	2	0	10uH
.TRAN 20us	50ms	0	20us
.PROBE
.END