PRACTICE_PROBLEM_3.CIR
I1	0	1	DC	2.0A
R1	1	0	2
R2	2	0	4
R3	1	2	10
V1	2	1	DC	2.0V
I2	2	0	DC	7.0A
.DC	V1	2	2	1
.PRINT	DC	V(1)	V(2)
.END
