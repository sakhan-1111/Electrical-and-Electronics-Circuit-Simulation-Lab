* C:\Users\Administrator\Desktop\Exam\3.sch

* Schematics Version 9.2
* Wed Dec 13 11:44:31 2017



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "3.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
