Lab_2_Ex_1.cir
R1	4	0	2
R2	2	3	3
R3	1	2	3
R4	1	3	10
E1	1	4	2	3	3
V1	3	0	DC 20V
I1 0	2	DC 0.1A
.DC V1 20 20 1
.PRINT DC V(2,3) I(E1)
.END