LAB-3-EXAMPLE-1-SOURCE.CIR
R1	1	3	5
R2	2	3	5
R3	2	0	10
R4	4	3	20
R5	3	5	10
RL 5	0	10
V1	1	0	DC	10V
I1	0	4	DC	1A
G1	0	3	2	0	2
.DC	LIN	V1	0	20	1
.PROBE
.END