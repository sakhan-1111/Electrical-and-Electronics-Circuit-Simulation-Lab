Practice_Problem_1.CIR
IDC4 0	63	DC	1.0A
R4	63	0	10
V7 63	67	DC 6.0V
R6	67	0	5
R8	67 68 7
V5 68 0 DC	2.0V
.DC V7 6	6	1	V5 2	2	1
.PRINT DC V(63) v(67) v(68)
.PRINT DC V(63,0)	I(R4)
.PRINT DC V(67,0)	I(R6)
.PRINT DC V(67,68) I(R8)
.END
