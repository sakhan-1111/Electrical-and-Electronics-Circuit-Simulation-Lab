Lab-5-Example-1-Netlist.cir
V1	1	0	DC	0	AC	0	SIN	0	100V	60Hz	0	0	0
C1	3	0	1uF
R1	1	2	1k
L1	2	3	10H
.TRAN 20us	50ms	0	20us
.PROBE
.END
