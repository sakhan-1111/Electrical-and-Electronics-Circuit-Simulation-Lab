Example_1.CIR 
Vs	1	0	DC	20.0V ; note the node placements 
Ra	1	2	5.0k
Rb	2	0	4.0k
Rc	3	0	1.0k
Is	3	2	DC	2.0mA ; note the node placements
.DC	Vs	20	20	1 ; this enables the .print commands
.PRINT	DC	V(1,2)	I(Ra)
.PRINT	DC	V(2)	I(Rb) 
.PRINT	DC	V(3)	I(Rc)
.END
