Lab_2_Exercise_2.cir
R1	1	2	8
R2	2	5	16
R3	6	0	4
R4	3	4	20
R5	4	0	8
V1	1	0	DC 10V
V2	5	6	DC 0V
F1	3	2	V2	0.5
.DC V1	10	10	1
.PRINT DC I(R2) V(3,2)
.END
