Lab_2_Example_3.cir
V1	1	0	DC 10
R1	1	2	8
R2	3	4	20
R3	0	4	8
R4	5	2	16
R5	0	5	4
F1	3	2	V1	0.5
.DC V1 10 10 1
.PRINT DC I(R1)
.END
