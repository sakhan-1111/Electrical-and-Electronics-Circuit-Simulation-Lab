Lab_4_Exercise_1_2.CIR
V1	1	0	DC	10V
R1	1	2	1k
Lag	2	0	1mH	IC=5mA
.TRAN	20us	0.02ms	0ms	10us	UIC
.PROBE
.END
