PRACTICE_PROBLEM_2.CIR
V1	1	0	DC 6.0V
R1	1	2	2
R4 1	3	4
R2	2	0	4
R3	2	3	6
I1 0	3	DC 4.0A
.DC V1 6 6 1
.PRINT DC V(1,2) I(R1)
.END
