EXANPLE-2-NETLIST.CIR
R1	0 1  1k 
I1	0 1 DC 10mA
C1	0 1  1uF IC=0V
.TRAN	20us	15ms	0ms	10us UIC
.PROBE
.END
